library verilog;
use verilog.vl_types.all;
entity ClkDiv_tb is
end ClkDiv_tb;
