module serializer #(parameter IN_WIDTH=8) (
input wire CLK,
input wire RST,
input wire [IN_WIDTH-1:0] P_DATA,
input wire DATA_VALID,
input wire ser_en,
input wire BUSY,
output reg ser_done,
output reg ser_data
);

integer j;
integer Counter ;
reg [IN_WIDTH-1:0] LFSR;
  

always@(posedge CLK or negedge RST)
begin
	if (!RST) 
		begin
			ser_data <= 1'b0;
			ser_done <= 1'b0;
			Counter<=0;
		end
		else if(DATA_VALID && !BUSY)
		  			begin
		  			LFSR <= P_DATA;
		  			end
		  			else if(ser_en && BUSY)
		begin
			 ser_data<= LFSR[0];  //Output takes the LSB
			
			//Loop on the register bits to shift right one bit
			for (j=0; j<=6; j=j+1)
			 LFSR [j] <= LFSR[j+1];    //High during the output operation
			if(Counter != 8)
			 Counter <= Counter+1;
			else
			  ser_done <= 1'b1;
	 	end
	else
		begin
			ser_data <= 1'b0;
			ser_done <= 1'b0;
			Counter<=0;
		end
					   
					       end
			     endmodule
		  
		  
		  
		

