module UART_TX(
input wire DATA_VALID,
input wire PAR_EN,
input wire ser_done,
input wire CLK,
input wire RST, 
output reg ser_en,
output reg BUSY,
output reg [1:0] mux_sel
);
localparam  [1:0]    IDLE = 2'b00,
                     START = 2'b01,
                     DATA = 2'b10,
                     PARITY=2'b11;
reg    [1:0]         current_state,
                     next_state ;
// state transition 		
always @(posedge CLK or negedge RST)
 begin
  if(!RST)
   begin
     current_state <= IDLE ;
   end
  else
   begin
     current_state <= next_state ;
   end
 end
 
// next_state logic
always @(*)
 begin
  case(current_state)
  IDLE     : begin
               if(DATA_VALID==1'b1&& ser_done==1'b0)
               begin
               next_state = START ;
               end	 
              else
			        next_state = IDLE ;         		  
             end
  START       :  next_state = DATA ;
	              
  DATA      : begin
              if(ser_done==1'b1&&PAR_EN==1'b0)
			          next_state = IDLE ;
			        else if(ser_done==1'b1&&PAR_EN==1'b1)
               next_state = PARITY ;
	              else
	                 next_state = DATA ;
	              end
	                
	 PARITY     : begin
                next_state = IDLE;
                end              
  default :   next_state = IDLE ;		 
  
  endcase
end	   
// output logic
always @(*)
 begin
   ser_en=1'b0;
   BUSY=1'b0;
   mux_sel=2'b01;
  case(current_state)
  IDLE     : begin
              if(DATA_VALID==1'b1)
                begin
              ser_en=1'b1;
              BUSY=1'b0;
               end
            else
              begin
              ser_en=1'b0; 
              BUSY=1'b0; 
              end
             end
  START       : begin
              mux_sel=2'b00;
              ser_en=1'b1;
              BUSY=1'b1;
               end
  DATA     : begin
               if(ser_done==1'b0)
               begin
                 mux_sel=2'b10;
                BUSY=1'b1;
                ser_en=1'b1;
               end
            else if(ser_done==1'b1&&PAR_EN==1'b0)
                begin
              mux_sel=2'b01;
              BUSY=1'b1;
              ser_en=1'b0;
              end
            else if(ser_done==1'b1&&PAR_EN==1'b1)
              begin
              mux_sel=2'b11; 
              BUSY=1'b1; 
              ser_en=1'b0;
             end 	   
             end
   PARITY     : begin
                mux_sel=2'b01;
                end
                
  default  : begin
              ser_en=1'b0;
              BUSY=1'b0;
              mux_sel=2'b01;
             end			  
  endcase
 end	
		
		
endmodule